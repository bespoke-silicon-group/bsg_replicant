`ifndef CL_TARGET_DEFINES
`define CL_TARGET_DEFINES

`define BSG_TARGET_F1

`endif
