// Amazon FPGA Hardware Development Kit
//
// Copyright 2016 Amazon.com, Inc. or its affiliates. All Rights Reserved.
//
// Licensed under the Amazon Software License (the "License"). You may not use
// this file except in compliance with the License. A copy of the License is
// located at
//
//    http://aws.amazon.com/asl/
//
// or in the "license" file accompanying this file. This file is distributed on
// an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, express or
// implied. See the License for the specific language governing permissions and
// limitations under the License.


module cl_fsb_tb();

import tb_type_defines_pkg::*;
`include "cl_common_defines.vh" // CL Defines with register addresses

// AXI ID
parameter [5:0] AXI_ID = 6'h0;

logic [31:0] rdata;
logic [15:0] vdip_value;
logic [15:0] vled_value;


   initial begin

      tb.power_up();
      #10 $display("Code modification");
      
      #10 tb.set_virtual_dip_switch(.dip(0));
      
      #10 vdip_value = tb.get_virtual_dip_switch();
      #10 $display ("value of vdip:%0x", vdip_value);
      $display ("Writing 0xDEAD_BEEF to address 0x%x", `DEMO_REG_ADDR);
      tb.poke(.addr(`DEMO_REG_ADDR), .data(32'hDEAD_BEEF), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL)); // write register
      # 10;
      tb.peek(.addr(`DEMO_REG_ADDR), .data(rdata), .id(AXI_ID), .size(DataSize::UINT16), .intf(AxiPort::PORT_OCL));         // start read & write
      $display ("Reading 0x%x from address 0x%x", rdata, `DEMO_REG_ADDR);
      # 10;
      if (rdata == 32'hEFBE_ADDE) // Check for byte swap in register read
        $display ("TEST PASSED");
      else
        $display ("TEST FAILED");
      # 10;
      tb.peek_ocl(.addr(`VLED_REG_ADDR), .data(rdata));         // start read
      $display ("Reading 0x%x from address 0x%x", rdata, `VLED_REG_ADDR);
      # 10;
      if (rdata == 32'h0000_BEEF) // Check for LED register read
        $display ("TEST PASSED");
      else
        $display ("TEST FAILED");
      # 10;
      vled_value = tb.get_virtual_led();
      # 10;
      $display ("value of vled:%0x", vled_value);

      tb.kernel_reset();
      # 10;
      tb.power_down();
      $display("%d", $stime);
      
      $finish;
   end

endmodule // test_cl_fsb
