/**
*  axi_perf_mon.v
*
*/

`include "bsg_axi_bus_pkg.vh"

module axi_perf_mon #(
  parameter slot_num_p = "inv"
  , parameter id_width_p = "inv"
  , parameter addr_width_p = "inv"
  , parameter data_width_p = "inv"
  , localparam axil_mosi_bus_width_lp = `bsg_axil_mosi_bus_width(1)
  , localparam axil_miso_bus_width_lp = `bsg_axil_miso_bus_width(1)
  , localparam axi_mosi_bus_width_lp = `bsg_axi_mosi_bus_width(1, id_width_p, addr_width_p, data_width_p)
  , localparam axi_miso_bus_width_lp = `bsg_axi_miso_bus_width(1, id_width_p, addr_width_p, data_width_p)
) (
  input                               s_axil_clk_i
  ,
  input                               s_axil_resetn_i
  ,
  input  [axil_mosi_bus_width_lp-1:0] s_axil_bus_i
  ,
  output [axil_miso_bus_width_lp-1:0] s_axil_bus_o
  ,
  input                               slot_0_axi_aclk_i
  ,
  input                               slot_0_axi_resetn_i
  ,
  input  [ axi_mosi_bus_width_lp-1:0] slot_0_axi_mo_i
  ,
  input  [ axi_miso_bus_width_lp-1:0] slot_0_axi_mi_i
  ,
  input                               core_clk_i
  ,
  input                               core_aresetn_i
  ,
  input                               capture_event_i
  ,
  input                               reset_event_i
  ,
  output                              interrupt_o
);


  `declare_bsg_axil_bus_s(1, bsg_s_axil_i_bus_s, bsg_s_axil_o_bus_s);
  bsg_s_axil_i_bus_s s_axil_bus_li_cast;
  bsg_s_axil_o_bus_s s_axil_bus_lo_cast;

  assign s_axil_bus_li_cast = s_axil_bus_i;
  assign s_axil_bus_o       = s_axil_bus_lo_cast;

  `declare_bsg_axi_bus_s(1, id_width_p, addr_width_p, data_width_p, bsg_axi_mosi_mux_s, bsg_axi_miso_mux_s);
  bsg_axi_mosi_mux_s axi_mo_cast;
  bsg_axi_miso_mux_s axi_mi_cast;

  assign axi_mo_cast = slot_0_axi_mo_i;
  assign axi_mi_cast = slot_0_axi_mi_i;

  axi_perf_mon_v5_0_19_top #(
    `ifdef BSG_TARGET_F1
    .C_FAMILY                    ("virtexuplus" ),
    `else
    .C_FAMILY                    ("virtexuplusHBM"),
    `endif
    .C_INSTANCE                  ("axi_perf_mon"),
    .C_LITE_ADDRESS_WIDTH        (16            ),
    .C_S_AXI_ADDR_WIDTH          (16            ),
    .C_S_AXI_DATA_WIDTH          (32            ),
    .C_S_AXI_PROTOCOL            ("AXI4LITE"    ),
    .C_S_AXI_ID_WIDTH            (1             ),
    .C_SUPPORT_ID_REFLECTION     (0             ),
    .C_ENABLE_ADVANCED           (1             ),
    .C_ENABLE_PROFILE            (0             ),
    .C_ENABLE_TRACE              (0             ),
    .C_EN_AXI_DEBUG              (0             ),
    .C_EN_TRIGGER                (0             ),
    .C_EN_WR_ADD_FLAG            (1             ),
    .C_EN_FIRST_WRITE_FLAG       (1             ),
    .C_EN_LAST_WRITE_FLAG        (1             ),
    .C_EN_RESPONSE_FLAG          (1             ),
    .C_EN_RD_ADD_FLAG            (1             ),
    .C_EN_FIRST_READ_FLAG        (1             ),
    .C_EN_LAST_READ_FLAG         (1             ),
    .C_EN_SW_REG_WR_FLAG         (0             ),
    .C_EN_EXT_EVENTS_FLAG        (0             ),
    .C_NUM_MONITOR_SLOTS         (slot_num_p    ),
    .C_ENABLE_EVENT_COUNT        (1             ),
    .C_NUM_OF_COUNTERS           (1             ),
    .C_METRIC_COUNT_WIDTH        (32            ),
    .C_METRIC_COUNT_SCALE        (1             ),
    .C_GLOBAL_COUNT_WIDTH        (64            ),
    .C_HAVE_SAMPLED_METRIC_CNT   (1             ),
    .C_METRICS_SAMPLE_COUNT_WIDTH(32            ),
    .C_AXI4LITE_CORE_CLK_ASYNC   (1             ),
    .C_SLOT_0_AXI_ADDR_WIDTH     (addr_width_p  ),
    .C_SLOT_0_AXI_DATA_WIDTH     (data_width_p  ),
    .C_SLOT_0_AXI_ID_WIDTH       (id_width_p    ),
    .C_SLOT_0_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_0_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_0_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_0_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_0_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_0_FIFO_ENABLE        (1             ),
    .C_SLOT_1_AXI_ADDR_WIDTH     (32            ),
    .C_SLOT_1_AXI_DATA_WIDTH     (32            ),
    .C_SLOT_1_AXI_ID_WIDTH       (1             ),
    .C_SLOT_1_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_1_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_1_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_1_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_1_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_1_FIFO_ENABLE        (1             ),
    .C_SLOT_2_AXI_ADDR_WIDTH     (32            ),
    .C_SLOT_2_AXI_DATA_WIDTH     (32            ),
    .C_SLOT_2_AXI_ID_WIDTH       (1             ),
    .C_SLOT_2_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_2_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_2_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_2_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_2_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_2_FIFO_ENABLE        (1             ),
    .C_SLOT_3_AXI_ADDR_WIDTH     (32            ),
    .C_SLOT_3_AXI_DATA_WIDTH     (32            ),
    .C_SLOT_3_AXI_ID_WIDTH       (1             ),
    .C_SLOT_3_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_3_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_3_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_3_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_3_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_3_FIFO_ENABLE        (1             ),
    .C_SLOT_4_AXI_ADDR_WIDTH     (32            ),
    .C_SLOT_4_AXI_DATA_WIDTH     (32            ),
    .C_SLOT_4_AXI_ID_WIDTH       (1             ),
    .C_SLOT_4_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_4_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_4_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_4_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_4_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_4_FIFO_ENABLE        (1             ),
    .C_SLOT_5_AXI_ADDR_WIDTH     (32            ),
    .C_SLOT_5_AXI_DATA_WIDTH     (32            ),
    .C_SLOT_5_AXI_ID_WIDTH       (1             ),
    .C_SLOT_5_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_5_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_5_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_5_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_5_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_5_FIFO_ENABLE        (1             ),
    .C_SLOT_6_AXI_ADDR_WIDTH     (32            ),
    .C_SLOT_6_AXI_DATA_WIDTH     (32            ),
    .C_SLOT_6_AXI_ID_WIDTH       (1             ),
    .C_SLOT_6_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_6_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_6_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_6_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_6_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_6_FIFO_ENABLE        (1             ),
    .C_SLOT_7_AXI_ADDR_WIDTH     (32            ),
    .C_SLOT_7_AXI_DATA_WIDTH     (32            ),
    .C_SLOT_7_AXI_ID_WIDTH       (1             ),
    .C_SLOT_7_AXI_PROTOCOL       ("AXI4"        ),
    .C_SLOT_7_AXIS_TDATA_WIDTH   (32            ),
    .C_SLOT_7_AXIS_TID_WIDTH     (1             ),
    .C_SLOT_7_AXIS_TDEST_WIDTH   (1             ),
    .C_SLOT_7_AXIS_TUSER_WIDTH   (1             ),
    .C_SLOT_7_FIFO_ENABLE        (1             ),
    .C_SLOT_0_AXI_AWLEN          (7             ),
    .C_SLOT_1_AXI_AWLEN          (7             ),
    .C_SLOT_2_AXI_AWLEN          (7             ),
    .C_SLOT_3_AXI_AWLEN          (7             ),
    .C_SLOT_4_AXI_AWLEN          (7             ),
    .C_SLOT_5_AXI_AWLEN          (7             ),
    .C_SLOT_6_AXI_AWLEN          (7             ),
    .C_SLOT_7_AXI_AWLEN          (7             ),
    .C_SLOT_0_AXI_LOCK           (0             ),
    .C_SLOT_1_AXI_LOCK           (0             ),
    .C_SLOT_2_AXI_LOCK           (0             ),
    .C_SLOT_3_AXI_LOCK           (0             ),
    .C_SLOT_4_AXI_LOCK           (0             ),
    .C_SLOT_5_AXI_LOCK           (0             ),
    .C_SLOT_6_AXI_LOCK           (0             ),
    .C_SLOT_7_AXI_LOCK           (0             ),
    .C_REG_ALL_MONITOR_SIGNALS   (0             ),
    .C_EXT_EVENT0_FIFO_ENABLE    (1             ),
    .C_EXT_EVENT1_FIFO_ENABLE    (1             ),
    .C_EXT_EVENT2_FIFO_ENABLE    (1             ),
    .C_EXT_EVENT3_FIFO_ENABLE    (1             ),
    .C_EXT_EVENT4_FIFO_ENABLE    (1             ),
    .C_EXT_EVENT5_FIFO_ENABLE    (1             ),
    .C_EXT_EVENT6_FIFO_ENABLE    (1             ),
    .C_EXT_EVENT7_FIFO_ENABLE    (1             ),
    .C_ENABLE_EVENT_LOG          (0             ),
    .C_FIFO_AXIS_DEPTH           (32            ),
    .C_FIFO_AXIS_TDATA_WIDTH     (56            ),
    .C_AXIS_DWIDTH_ROUND_TO_32   (64            ),
    .C_FIFO_AXIS_TID_WIDTH       (1             ),
    .C_FIFO_AXIS_SYNC            (0             ),
    .C_SHOW_AXI_IDS              (0             ),
    .C_SHOW_AXI_LEN              (0             ),
    .C_SHOW_AXIS_TID             (0             ),
    .C_SHOW_AXIS_TDEST           (0             ),
    .C_SHOW_AXIS_TUSER           (0             ),
    .ENABLE_EXT_EVENTS           (0             ),
    .COUNTER_LOAD_VALUE          ('H00000000    ),
    .C_LOG_DATA_OFFLD            (0             ),
    .S_AXI_OFFLD_ID_WIDTH        (1             ),
    .C_S_AXI4_BASEADDR           ('HFFFFFFFF    ),
    .C_S_AXI4_HIGHADDR           ('H00000000    ),
    .C_EN_ALL_TRACE              (1             )
  ) axi_perf_mon (
    .s_axi_aclk           (s_axil_clk_i                   ),
    .s_axi_aresetn        (s_axil_resetn_i                ),
    .s_axi_awaddr         (s_axil_bus_li_cast.awaddr[15:0]),
    .s_axi_awvalid        (s_axil_bus_li_cast.awvalid     ),
    .s_axi_awid           (1'B0                           ),
    .s_axi_awready        (s_axil_bus_lo_cast.awready     ),
    .s_axi_wdata          (s_axil_bus_li_cast.wdata       ),
    .s_axi_wstrb          (s_axil_bus_li_cast.wstrb       ),
    .s_axi_wvalid         (s_axil_bus_li_cast.wvalid      ),
    .s_axi_wready         (s_axil_bus_lo_cast.wready      ),
    .s_axi_bresp          (s_axil_bus_lo_cast.bresp       ),
    .s_axi_bvalid         (s_axil_bus_lo_cast.bvalid      ),
    .s_axi_bid            (                               ),
    .s_axi_bready         (s_axil_bus_li_cast.bready      ),
    .s_axi_araddr         (s_axil_bus_li_cast.araddr[15:0]),
    .s_axi_arvalid        (s_axil_bus_li_cast.arvalid     ),
    .s_axi_arid           (1'B0                           ),
    .s_axi_arready        (s_axil_bus_lo_cast.arready     ),
    .s_axi_rdata          (s_axil_bus_lo_cast.rdata       ),
    .s_axi_rresp          (s_axil_bus_lo_cast.rresp       ),
    .s_axi_rvalid         (s_axil_bus_lo_cast.rvalid      ),
    .s_axi_rid            (                               ),
    .s_axi_rready         (s_axil_bus_li_cast.rready      ),
    
    .slot_0_axi_aclk      (slot_0_axi_aclk_i              ),
    .slot_0_axi_aresetn   (slot_0_axi_resetn_i            ),
    .slot_0_axi_awid      (axi_mo_cast.awid               ),
    .slot_0_axi_awaddr    (axi_mo_cast.awaddr             ),
    .slot_0_axi_awprot    (axi_mo_cast.awprot             ),
    .slot_0_axi_awlen     (axi_mo_cast.awlen              ),
    .slot_0_axi_awsize    (axi_mo_cast.awsize             ),
    .slot_0_axi_awburst   (axi_mo_cast.awburst            ),
    .slot_0_axi_awcache   (axi_mo_cast.awcache            ),
    .slot_0_axi_awlock    (axi_mo_cast.awlock             ),
    .slot_0_axi_awvalid   (axi_mo_cast.awvalid            ),
    .slot_0_axi_awready   (axi_mi_cast.awready            ),
    .slot_0_axi_wdata     (axi_mo_cast.wdata              ),
    .slot_0_axi_wstrb     (axi_mo_cast.wstrb              ),
    .slot_0_axi_wlast     (axi_mo_cast.wlast              ),
    .slot_0_axi_wvalid    (axi_mo_cast.wvalid             ),
    .slot_0_axi_wready    (axi_mi_cast.wready             ),
    .slot_0_axi_bid       (axi_mi_cast.bid                ),
    .slot_0_axi_bresp     (axi_mi_cast.bresp              ),
    .slot_0_axi_bvalid    (axi_mi_cast.bvalid             ),
    .slot_0_axi_bready    (axi_mo_cast.bready             ),
    .slot_0_axi_arid      (axi_mo_cast.arid               ),
    .slot_0_axi_araddr    (axi_mo_cast.araddr             ),
    .slot_0_axi_arlen     (axi_mo_cast.arlen              ),
    .slot_0_axi_arsize    (axi_mo_cast.arsize             ),
    .slot_0_axi_arburst   (axi_mo_cast.arburst            ),
    .slot_0_axi_arcache   (axi_mo_cast.arcache            ),
    .slot_0_axi_arprot    (axi_mo_cast.arprot             ),
    .slot_0_axi_arlock    (axi_mo_cast.arlock             ),
    .slot_0_axi_arvalid   (axi_mo_cast.arvalid            ),
    .slot_0_axi_arready   (axi_mi_cast.arready            ),
    .slot_0_axi_rid       (axi_mi_cast.rid                ),
    .slot_0_axi_rdata     (axi_mi_cast.rdata              ),
    .slot_0_axi_rresp     (axi_mi_cast.rresp              ),
    .slot_0_axi_rlast     (axi_mi_cast.rlast              ),
    .slot_0_axi_rvalid    (axi_mi_cast.rvalid             ),
    .slot_0_axi_rready    (axi_mo_cast.rready             ),
    .slot_0_axis_aclk     (1'B0                           ),
    .slot_0_axis_aresetn  (1'B1                           ),
    .slot_0_axis_tvalid   (1'B0                           ),
    .slot_0_axis_tready   (1'B0                           ),
    .slot_0_axis_tdata    (32'B0                          ),
    .slot_0_axis_tstrb    (4'HF                           ),
    .slot_0_axis_tkeep    (4'HF                           ),
    .slot_0_axis_tlast    (1'B0                           ),
    .slot_0_axis_tid      (1'B0                           ),
    .slot_0_axis_tdest    (1'B0                           ),
    .slot_0_axis_tuser    (1'B0                           ),
    .slot_0_ext_trig      (1'B0                           ),
    .slot_0_ext_trig_stop (1'B0                           ),
    
    .slot_1_axi_aclk      (1'B0                           ),
    .slot_1_axi_aresetn   (1'B1                           ),
    .slot_1_axi_awid      (1'B0                           ),
    .slot_1_axi_awaddr    (32'B0                          ),
    .slot_1_axi_awprot    (3'B0                           ),
    .slot_1_axi_awlen     (8'B0                           ),
    .slot_1_axi_awsize    (3'B0                           ),
    .slot_1_axi_awburst   (2'B0                           ),
    .slot_1_axi_awcache   (4'B0                           ),
    .slot_1_axi_awlock    (1'B0                           ),
    .slot_1_axi_awvalid   (1'B0                           ),
    .slot_1_axi_awready   (1'B0                           ),
    .slot_1_axi_wdata     (32'B0                          ),
    .slot_1_axi_wstrb     (4'B0                           ),
    .slot_1_axi_wlast     (1'B0                           ),
    .slot_1_axi_wvalid    (1'B0                           ),
    .slot_1_axi_wready    (1'B0                           ),
    .slot_1_axi_bid       (1'B0                           ),
    .slot_1_axi_bresp     (2'B0                           ),
    .slot_1_axi_bvalid    (1'B0                           ),
    .slot_1_axi_bready    (1'B0                           ),
    .slot_1_axi_arid      (1'B0                           ),
    .slot_1_axi_araddr    (32'B0                          ),
    .slot_1_axi_arlen     (8'B0                           ),
    .slot_1_axi_arsize    (3'B0                           ),
    .slot_1_axi_arburst   (2'B0                           ),
    .slot_1_axi_arcache   (4'B0                           ),
    .slot_1_axi_arprot    (3'B0                           ),
    .slot_1_axi_arlock    (1'B0                           ),
    .slot_1_axi_arvalid   (1'B0                           ),
    .slot_1_axi_arready   (1'B0                           ),
    .slot_1_axi_rid       (1'B0                           ),
    .slot_1_axi_rdata     (32'B0                          ),
    .slot_1_axi_rresp     (2'B0                           ),
    .slot_1_axi_rlast     (1'B0                           ),
    .slot_1_axi_rvalid    (1'B0                           ),
    .slot_1_axi_rready    (1'B0                           ),
    .slot_1_axis_aclk     (1'B0                           ),
    .slot_1_axis_aresetn  (1'B1                           ),
    .slot_1_axis_tvalid   (1'B0                           ),
    .slot_1_axis_tready   (1'B0                           ),
    .slot_1_axis_tdata    (32'B0                          ),
    .slot_1_axis_tstrb    (4'HF                           ),
    .slot_1_axis_tkeep    (4'HF                           ),
    .slot_1_axis_tlast    (1'B0                           ),
    .slot_1_axis_tid      (1'B0                           ),
    .slot_1_axis_tdest    (1'B0                           ),
    .slot_1_axis_tuser    (1'B0                           ),
    .slot_1_ext_trig      (1'B0                           ),
    .slot_1_ext_trig_stop (1'B0                           ),
    .slot_2_axi_aclk      (1'B0                           ),
    .slot_2_axi_aresetn   (1'B1                           ),
    .slot_2_axi_awid      (1'B0                           ),
    .slot_2_axi_awaddr    (32'B0                          ),
    .slot_2_axi_awprot    (3'B0                           ),
    .slot_2_axi_awlen     (8'B0                           ),
    .slot_2_axi_awsize    (3'B0                           ),
    .slot_2_axi_awburst   (2'B0                           ),
    .slot_2_axi_awcache   (4'B0                           ),
    .slot_2_axi_awlock    (1'B0                           ),
    .slot_2_axi_awvalid   (1'B0                           ),
    .slot_2_axi_awready   (1'B0                           ),
    .slot_2_axi_wdata     (32'B0                          ),
    .slot_2_axi_wstrb     (4'B0                           ),
    .slot_2_axi_wlast     (1'B0                           ),
    .slot_2_axi_wvalid    (1'B0                           ),
    .slot_2_axi_wready    (1'B0                           ),
    .slot_2_axi_bid       (1'B0                           ),
    .slot_2_axi_bresp     (2'B0                           ),
    .slot_2_axi_bvalid    (1'B0                           ),
    .slot_2_axi_bready    (1'B0                           ),
    .slot_2_axi_arid      (1'B0                           ),
    .slot_2_axi_araddr    (32'B0                          ),
    .slot_2_axi_arlen     (8'B0                           ),
    .slot_2_axi_arsize    (3'B0                           ),
    .slot_2_axi_arburst   (2'B0                           ),
    .slot_2_axi_arcache   (4'B0                           ),
    .slot_2_axi_arprot    (3'B0                           ),
    .slot_2_axi_arlock    (1'B0                           ),
    .slot_2_axi_arvalid   (1'B0                           ),
    .slot_2_axi_arready   (1'B0                           ),
    .slot_2_axi_rid       (1'B0                           ),
    .slot_2_axi_rdata     (32'B0                          ),
    .slot_2_axi_rresp     (2'B0                           ),
    .slot_2_axi_rlast     (1'B0                           ),
    .slot_2_axi_rvalid    (1'B0                           ),
    .slot_2_axi_rready    (1'B0                           ),
    .slot_2_axis_aclk     (1'B0                           ),
    .slot_2_axis_aresetn  (1'B1                           ),
    .slot_2_axis_tvalid   (1'B0                           ),
    .slot_2_axis_tready   (1'B0                           ),
    .slot_2_axis_tdata    (32'B0                          ),
    .slot_2_axis_tstrb    (4'HF                           ),
    .slot_2_axis_tkeep    (4'HF                           ),
    .slot_2_axis_tlast    (1'B0                           ),
    .slot_2_axis_tid      (1'B0                           ),
    .slot_2_axis_tdest    (1'B0                           ),
    .slot_2_axis_tuser    (1'B0                           ),
    .slot_2_ext_trig      (1'B0                           ),
    .slot_2_ext_trig_stop (1'B0                           ),
    .slot_3_axi_aclk      (1'B0                           ),
    .slot_3_axi_aresetn   (1'B1                           ),
    .slot_3_axi_awid      (1'B0                           ),
    .slot_3_axi_awaddr    (32'B0                          ),
    .slot_3_axi_awprot    (3'B0                           ),
    .slot_3_axi_awlen     (8'B0                           ),
    .slot_3_axi_awsize    (3'B0                           ),
    .slot_3_axi_awburst   (2'B0                           ),
    .slot_3_axi_awcache   (4'B0                           ),
    .slot_3_axi_awlock    (1'B0                           ),
    .slot_3_axi_awvalid   (1'B0                           ),
    .slot_3_axi_awready   (1'B0                           ),
    .slot_3_axi_wdata     (32'B0                          ),
    .slot_3_axi_wstrb     (4'B0                           ),
    .slot_3_axi_wlast     (1'B0                           ),
    .slot_3_axi_wvalid    (1'B0                           ),
    .slot_3_axi_wready    (1'B0                           ),
    .slot_3_axi_bid       (1'B0                           ),
    .slot_3_axi_bresp     (2'B0                           ),
    .slot_3_axi_bvalid    (1'B0                           ),
    .slot_3_axi_bready    (1'B0                           ),
    .slot_3_axi_arid      (1'B0                           ),
    .slot_3_axi_araddr    (32'B0                          ),
    .slot_3_axi_arlen     (8'B0                           ),
    .slot_3_axi_arsize    (3'B0                           ),
    .slot_3_axi_arburst   (2'B0                           ),
    .slot_3_axi_arcache   (4'B0                           ),
    .slot_3_axi_arprot    (3'B0                           ),
    .slot_3_axi_arlock    (1'B0                           ),
    .slot_3_axi_arvalid   (1'B0                           ),
    .slot_3_axi_arready   (1'B0                           ),
    .slot_3_axi_rid       (1'B0                           ),
    .slot_3_axi_rdata     (32'B0                          ),
    .slot_3_axi_rresp     (2'B0                           ),
    .slot_3_axi_rlast     (1'B0                           ),
    .slot_3_axi_rvalid    (1'B0                           ),
    .slot_3_axi_rready    (1'B0                           ),
    .slot_3_axis_aclk     (1'B0                           ),
    .slot_3_axis_aresetn  (1'B1                           ),
    .slot_3_axis_tvalid   (1'B0                           ),
    .slot_3_axis_tready   (1'B0                           ),
    .slot_3_axis_tdata    (32'B0                          ),
    .slot_3_axis_tstrb    (4'HF                           ),
    .slot_3_axis_tkeep    (4'HF                           ),
    .slot_3_axis_tlast    (1'B0                           ),
    .slot_3_axis_tid      (1'B0                           ),
    .slot_3_axis_tdest    (1'B0                           ),
    .slot_3_axis_tuser    (1'B0                           ),
    .slot_3_ext_trig      (1'B0                           ),
    .slot_3_ext_trig_stop (1'B0                           ),
    .slot_4_axi_aclk      (1'B0                           ),
    .slot_4_axi_aresetn   (1'B1                           ),
    .slot_4_axi_awid      (1'B0                           ),
    .slot_4_axi_awaddr    (32'B0                          ),
    .slot_4_axi_awprot    (3'B0                           ),
    .slot_4_axi_awlen     (8'B0                           ),
    .slot_4_axi_awsize    (3'B0                           ),
    .slot_4_axi_awburst   (2'B0                           ),
    .slot_4_axi_awcache   (4'B0                           ),
    .slot_4_axi_awlock    (1'B0                           ),
    .slot_4_axi_awvalid   (1'B0                           ),
    .slot_4_axi_awready   (1'B0                           ),
    .slot_4_axi_wdata     (32'B0                          ),
    .slot_4_axi_wstrb     (4'B0                           ),
    .slot_4_axi_wlast     (1'B0                           ),
    .slot_4_axi_wvalid    (1'B0                           ),
    .slot_4_axi_wready    (1'B0                           ),
    .slot_4_axi_bid       (1'B0                           ),
    .slot_4_axi_bresp     (2'B0                           ),
    .slot_4_axi_bvalid    (1'B0                           ),
    .slot_4_axi_bready    (1'B0                           ),
    .slot_4_axi_arid      (1'B0                           ),
    .slot_4_axi_araddr    (32'B0                          ),
    .slot_4_axi_arlen     (8'B0                           ),
    .slot_4_axi_arsize    (3'B0                           ),
    .slot_4_axi_arburst   (2'B0                           ),
    .slot_4_axi_arcache   (4'B0                           ),
    .slot_4_axi_arprot    (3'B0                           ),
    .slot_4_axi_arlock    (1'B0                           ),
    .slot_4_axi_arvalid   (1'B0                           ),
    .slot_4_axi_arready   (1'B0                           ),
    .slot_4_axi_rid       (1'B0                           ),
    .slot_4_axi_rdata     (32'B0                          ),
    .slot_4_axi_rresp     (2'B0                           ),
    .slot_4_axi_rlast     (1'B0                           ),
    .slot_4_axi_rvalid    (1'B0                           ),
    .slot_4_axi_rready    (1'B0                           ),
    .slot_4_axis_aclk     (1'B0                           ),
    .slot_4_axis_aresetn  (1'B1                           ),
    .slot_4_axis_tvalid   (1'B0                           ),
    .slot_4_axis_tready   (1'B0                           ),
    .slot_4_axis_tdata    (32'B0                          ),
    .slot_4_axis_tstrb    (4'HF                           ),
    .slot_4_axis_tkeep    (4'HF                           ),
    .slot_4_axis_tlast    (1'B0                           ),
    .slot_4_axis_tid      (1'B0                           ),
    .slot_4_axis_tdest    (1'B0                           ),
    .slot_4_axis_tuser    (1'B0                           ),
    .slot_4_ext_trig      (1'B0                           ),
    .slot_4_ext_trig_stop (1'B0                           ),
    .slot_5_axi_aclk      (1'B0                           ),
    .slot_5_axi_aresetn   (1'B0                           ),
    .slot_5_axi_awid      (1'B0                           ),
    .slot_5_axi_awaddr    (32'B0                          ),
    .slot_5_axi_awprot    (3'B0                           ),
    .slot_5_axi_awlen     (8'B0                           ),
    .slot_5_axi_awsize    (3'B0                           ),
    .slot_5_axi_awburst   (2'B0                           ),
    .slot_5_axi_awcache   (4'B0                           ),
    .slot_5_axi_awlock    (1'B0                           ),
    .slot_5_axi_awvalid   (1'B0                           ),
    .slot_5_axi_awready   (1'B0                           ),
    .slot_5_axi_wdata     (32'B0                          ),
    .slot_5_axi_wstrb     (4'B0                           ),
    .slot_5_axi_wlast     (1'B0                           ),
    .slot_5_axi_wvalid    (1'B0                           ),
    .slot_5_axi_wready    (1'B0                           ),
    .slot_5_axi_bid       (1'B0                           ),
    .slot_5_axi_bresp     (2'B0                           ),
    .slot_5_axi_bvalid    (1'B0                           ),
    .slot_5_axi_bready    (1'B0                           ),
    .slot_5_axi_arid      (1'B0                           ),
    .slot_5_axi_araddr    (32'B0                          ),
    .slot_5_axi_arlen     (8'B0                           ),
    .slot_5_axi_arsize    (3'B0                           ),
    .slot_5_axi_arburst   (2'B0                           ),
    .slot_5_axi_arcache   (4'B0                           ),
    .slot_5_axi_arprot    (3'B0                           ),
    .slot_5_axi_arlock    (1'B0                           ),
    .slot_5_axi_arvalid   (1'B0                           ),
    .slot_5_axi_arready   (1'B0                           ),
    .slot_5_axi_rid       (1'B0                           ),
    .slot_5_axi_rdata     (32'B0                          ),
    .slot_5_axi_rresp     (2'B0                           ),
    .slot_5_axi_rlast     (1'B0                           ),
    .slot_5_axi_rvalid    (1'B0                           ),
    .slot_5_axi_rready    (1'B0                           ),
    .slot_5_axis_aclk     (1'B0                           ),
    .slot_5_axis_aresetn  (1'B1                           ),
    .slot_5_axis_tvalid   (1'B0                           ),
    .slot_5_axis_tready   (1'B0                           ),
    .slot_5_axis_tdata    (32'B0                          ),
    .slot_5_axis_tstrb    (4'HF                           ),
    .slot_5_axis_tkeep    (4'HF                           ),
    .slot_5_axis_tlast    (1'B0                           ),
    .slot_5_axis_tid      (1'B0                           ),
    .slot_5_axis_tdest    (1'B0                           ),
    .slot_5_axis_tuser    (1'B0                           ),
    .slot_5_ext_trig      (1'B0                           ),
    .slot_5_ext_trig_stop (1'B0                           ),
    .slot_6_axi_aclk      (1'B0                           ),
    .slot_6_axi_aresetn   (1'B1                           ),
    .slot_6_axi_awid      (1'B0                           ),
    .slot_6_axi_awaddr    (32'B0                          ),
    .slot_6_axi_awprot    (3'B0                           ),
    .slot_6_axi_awlen     (8'B0                           ),
    .slot_6_axi_awsize    (3'B0                           ),
    .slot_6_axi_awburst   (2'B0                           ),
    .slot_6_axi_awcache   (4'B0                           ),
    .slot_6_axi_awlock    (1'B0                           ),
    .slot_6_axi_awvalid   (1'B0                           ),
    .slot_6_axi_awready   (1'B0                           ),
    .slot_6_axi_wdata     (32'B0                          ),
    .slot_6_axi_wstrb     (4'B0                           ),
    .slot_6_axi_wlast     (1'B0                           ),
    .slot_6_axi_wvalid    (1'B0                           ),
    .slot_6_axi_wready    (1'B0                           ),
    .slot_6_axi_bid       (1'B0                           ),
    .slot_6_axi_bresp     (2'B0                           ),
    .slot_6_axi_bvalid    (1'B0                           ),
    .slot_6_axi_bready    (1'B0                           ),
    .slot_6_axi_arid      (1'B0                           ),
    .slot_6_axi_araddr    (32'B0                          ),
    .slot_6_axi_arlen     (8'B0                           ),
    .slot_6_axi_arsize    (3'B0                           ),
    .slot_6_axi_arburst   (2'B0                           ),
    .slot_6_axi_arcache   (4'B0                           ),
    .slot_6_axi_arprot    (3'B0                           ),
    .slot_6_axi_arlock    (1'B0                           ),
    .slot_6_axi_arvalid   (1'B0                           ),
    .slot_6_axi_arready   (1'B0                           ),
    .slot_6_axi_rid       (1'B0                           ),
    .slot_6_axi_rdata     (32'B0                          ),
    .slot_6_axi_rresp     (2'B0                           ),
    .slot_6_axi_rlast     (1'B0                           ),
    .slot_6_axi_rvalid    (1'B0                           ),
    .slot_6_axi_rready    (1'B0                           ),
    .slot_6_axis_aclk     (1'B0                           ),
    .slot_6_axis_aresetn  (1'B1                           ),
    .slot_6_axis_tvalid   (1'B0                           ),
    .slot_6_axis_tready   (1'B0                           ),
    .slot_6_axis_tdata    (32'B0                          ),
    .slot_6_axis_tstrb    (4'HF                           ),
    .slot_6_axis_tkeep    (4'HF                           ),
    .slot_6_axis_tlast    (1'B0                           ),
    .slot_6_axis_tid      (1'B0                           ),
    .slot_6_axis_tdest    (1'B0                           ),
    .slot_6_axis_tuser    (1'B0                           ),
    .slot_6_ext_trig      (1'B0                           ),
    .slot_6_ext_trig_stop (1'B0                           ),
    .slot_7_axi_aclk      (1'B0                           ),
    .slot_7_axi_aresetn   (1'B1                           ),
    .slot_7_axi_awid      (1'B0                           ),
    .slot_7_axi_awaddr    (32'B0                          ),
    .slot_7_axi_awprot    (3'B0                           ),
    .slot_7_axi_awlen     (8'B0                           ),
    .slot_7_axi_awsize    (3'B0                           ),
    .slot_7_axi_awburst   (2'B0                           ),
    .slot_7_axi_awcache   (4'B0                           ),
    .slot_7_axi_awlock    (1'B0                           ),
    .slot_7_axi_awvalid   (1'B0                           ),
    .slot_7_axi_awready   (1'B0                           ),
    .slot_7_axi_wdata     (32'B0                          ),
    .slot_7_axi_wstrb     (4'B0                           ),
    .slot_7_axi_wlast     (1'B0                           ),
    .slot_7_axi_wvalid    (1'B0                           ),
    .slot_7_axi_wready    (1'B0                           ),
    .slot_7_axi_bid       (1'B0                           ),
    .slot_7_axi_bresp     (2'B0                           ),
    .slot_7_axi_bvalid    (1'B0                           ),
    .slot_7_axi_bready    (1'B0                           ),
    .slot_7_axi_arid      (1'B0                           ),
    .slot_7_axi_araddr    (32'B0                          ),
    .slot_7_axi_arlen     (8'B0                           ),
    .slot_7_axi_arsize    (3'B0                           ),
    .slot_7_axi_arburst   (2'B0                           ),
    .slot_7_axi_arcache   (4'B0                           ),
    .slot_7_axi_arprot    (3'B0                           ),
    .slot_7_axi_arlock    (1'B0                           ),
    .slot_7_axi_arvalid   (1'B0                           ),
    .slot_7_axi_arready   (1'B0                           ),
    .slot_7_axi_rid       (1'B0                           ),
    .slot_7_axi_rdata     (32'B0                          ),
    .slot_7_axi_rresp     (2'B0                           ),
    .slot_7_axi_rlast     (1'B0                           ),
    .slot_7_axi_rvalid    (1'B0                           ),
    .slot_7_axi_rready    (1'B0                           ),
    .slot_7_axis_aclk     (1'B0                           ),
    .slot_7_axis_aresetn  (1'B1                           ),
    .slot_7_axis_tvalid   (1'B0                           ),
    .slot_7_axis_tready   (1'B0                           ),
    .slot_7_axis_tdata    (32'B0                          ),
    .slot_7_axis_tstrb    (4'HF                           ),
    .slot_7_axis_tkeep    (4'HF                           ),
    .slot_7_axis_tlast    (1'B0                           ),
    .slot_7_axis_tid      (1'B0                           ),
    .slot_7_axis_tdest    (1'B0                           ),
    .slot_7_axis_tuser    (1'B0                           ),
    .slot_7_ext_trig      (1'B0                           ),
    .slot_7_ext_trig_stop (1'B0                           ),
    .ext_clk_0            (1'B0                           ),
    .ext_rstn_0           (1'B1                           ),
    .ext_event_0_cnt_start(1'B0                           ),
    .ext_event_0_cnt_stop (1'B0                           ),
    .ext_event_0          (1'B0                           ),
    .ext_clk_1            (1'B0                           ),
    .ext_rstn_1           (1'B1                           ),
    .ext_event_1_cnt_start(1'B0                           ),
    .ext_event_1_cnt_stop (1'B0                           ),
    .ext_event_1          (1'B0                           ),
    .ext_clk_2            (1'B0                           ),
    .ext_rstn_2           (1'B1                           ),
    .ext_event_2_cnt_start(1'B0                           ),
    .ext_event_2_cnt_stop (1'B0                           ),
    .ext_event_2          (1'B0                           ),
    .ext_clk_3            (1'B0                           ),
    .ext_rstn_3           (1'B1                           ),
    .ext_event_3_cnt_start(1'B0                           ),
    .ext_event_3_cnt_stop (1'B0                           ),
    .ext_event_3          (1'B0                           ),
    .ext_clk_4            (1'B0                           ),
    .ext_rstn_4           (1'B1                           ),
    .ext_event_4_cnt_start(1'B0                           ),
    .ext_event_4_cnt_stop (1'B0                           ),
    .ext_event_4          (1'B0                           ),
    .ext_clk_5            (1'B0                           ),
    .ext_rstn_5           (1'B1                           ),
    .ext_event_5_cnt_start(1'B0                           ),
    .ext_event_5_cnt_stop (1'B0                           ),
    .ext_event_5          (1'B0                           ),
    .ext_clk_6            (1'B0                           ),
    .ext_rstn_6           (1'B1                           ),
    .ext_event_6_cnt_start(1'B0                           ),
    .ext_event_6_cnt_stop (1'B0                           ),
    .ext_event_6          (1'B0                           ),
    .ext_clk_7            (1'B0                           ),
    .ext_rstn_7           (1'B1                           ),
    .ext_event_7_cnt_start(1'B0                           ),
    .ext_event_7_cnt_stop (1'B0                           ),
    .ext_event_7          (1'B0                           ),
    .capture_event        (capture_event_i                ),
    .reset_event          (reset_event_i                  ),
    .core_aclk            (core_clk_i                     ),
    .core_aresetn         (core_aresetn_i                 ),
    .m_axis_aclk          (1'B0                           ),
    .m_axis_aresetn       (1'B1                           ),
    .m_axis_tdata         (                               ),
    .m_axis_tstrb         (                               ),
    .m_axis_tvalid        (                               ),
    .m_axis_tid           (                               ),
    .m_axis_tready        (1'B0                           ),
    .s_axi_offld_aclk     (1'B0                           ),
    .s_axi_offld_aresetn  (1'B1                           ),
    .s_axi_offld_araddr   (32'B0                          ),
    .s_axi_offld_arvalid  (1'B0                           ),
    .s_axi_offld_arlen    (8'B0                           ),
    .s_axi_offld_arid     (1'B0                           ),
    .s_axi_offld_arready  (                               ),
    .s_axi_offld_rready   (1'B0                           ),
    .s_axi_offld_rdata    (                               ),
    .s_axi_offld_rresp    (                               ),
    .s_axi_offld_rvalid   (                               ),
    .s_axi_offld_rid      (                               ),
    .s_axi_offld_rlast    (                               ),
    .interrupt            (interrupt_o                    ),
    .trigger_in           (1'B0                           ),
    .trigger_in_ack       (                               )
  );

endmodule
